module test (
  // clock
  input clk,
  // reset
  input rst_n,
  // data
  input [63:0] d,
  output [63:0] q
);

endmodule
