module test (
);

endmodule
